module greater_than (
    A, B, F
);

input [1]
    
endmodule