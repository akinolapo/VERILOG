module greater_than (
    A, B, F
);
    
endmodule