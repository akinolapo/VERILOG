//2-to-4 Line Decoder
//4 AND gates on the output
//2x 1-to-2 Line Decoders

module moduleName (
    ports
);
    
endmodule