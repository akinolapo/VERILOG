module gre (
    ports
);
    
endmodule