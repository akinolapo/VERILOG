`timescale 1ns/1ns
`include "decoder.v"

module decoder1to2_tb;

reg A;
wire ;

endmodule