module hello (
    A, B
);

    input A
    
endmodule