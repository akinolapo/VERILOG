module hello (
    ports
);
    
endmodule