module greater_than (
    A, B, F
);

input []
    
endmodule