module hello (
    A, B
);

    input
    
endmodule