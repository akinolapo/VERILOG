module greater_than (
    A, B, C
);
    
endmodule