`timescale 1ns/1ns
`include "decoder.v"

module decoder2to4_tb;



endmodule