`timescale 1ps/1ps
`include "hello.v"

module hello_tb;