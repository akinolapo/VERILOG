module greater_than (
    A, B, F
);

in
    
endmodule