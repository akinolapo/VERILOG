module greater_than (
    A, B, F
);

input [1:0] A, B;
output F;

ass
    
endmodule