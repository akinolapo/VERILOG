module greater_than (
    ports
);
    
endmodule