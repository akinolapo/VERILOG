module hello (
    A, B
);

    input A;
    output B;
    
    
endmodule