module hello (
    A, B
);

    
    
endmodule