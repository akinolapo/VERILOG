module greater (
    ports
);
    
endmodule