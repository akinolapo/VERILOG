module hello (
    A, B
);

    inpu
    
endmodule