module hello (
    A, B
);

    input A;
    output B;

    assign
    
endmodule