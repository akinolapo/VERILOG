`timescale 1ps/1ps
`include "greater_than.v"

module greater_than_tb;

reg[1:0]
endmodule